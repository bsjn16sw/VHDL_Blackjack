library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity player is
end player;

architecture Behavioral of player is

begin


end Behavioral;

