library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity game is
end game;

architecture Behavioral of game is

begin


end Behavioral;

