library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity round is
end round;

architecture Behavioral of round is

begin


end Behavioral;

